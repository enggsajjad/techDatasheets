//*********************************************************************************************//
//    Project      : NexTek Service
//    File         : Uat_top.v
//    Author       : NexTek Service
//    Company      : NexTek Service
//    Start Date   : Nov  06th, 2004.
//    Last Updated : Dec  15th, 2004.
//    Version      : 2.0
//    Device	   : xc2s150-5pq208 
//    PROM	   : xcf01s
//    Abstract     : This is top level Module that defines Transmitter
// 
//    Modification History:
//==============================================================================================
//    Date                       By                 Version                Change Description
//==============================================================================================
//    Jan 01th, 2004          NexTek Service         0.1                   Original Version
//*********************************************************************************************//
 
// Desighn Block
module uat_top(//Inputs
               clk,                      //1-bit System Clock input
               rst_n,                    //1-bit Asyncronous Active Low Reset input
               din_rdy,                  //1-bit ready input signal that indicates the data is ready at input for Tx 
               din_byte,                 //8-bit data input in UART for Tx
               // Output
               ser_out,                  //1-bit Tx data output from UART
               uart_ready                //1-bit control signal goes to Sequence Controller                 
              );

// Declaration inputs, outputs 
input       clk;
input       rst_n;
input       din_rdy;
input [7:0] din_byte;    


output      ser_out;      
output      uart_ready;

reg         ser_out;

reg   [7:0] data_buf;         
reg   [2:0] shift_count;
reg         din_rdy_reg;
reg   [4:0] count ;
wire        start_bit_sig;
wire        data_bits_sig;
wire        stop_bit_sig;
      
// Registered Data Ready Signal
always @(negedge clk or negedge rst_n)
begin
  if(~rst_n)
    din_rdy_reg <= 1'b0;
  else
    din_rdy_reg <= din_rdy ; 
end 


//Output Logic
always @(negedge clk or negedge rst_n)
begin
   if(~rst_n)
      ser_out <= 1'b1;
   else 
   begin
     case({start_bit_sig,data_bits_sig,stop_bit_sig})
        3'b100: ser_out <= 1'b0;
        3'b010: ser_out <= data_buf[0];
        3'b001: ser_out <= 1'b1;
        default: ser_out <= 1'b1;
     endcase
   end
end         

// strat bit pipelinin
always @(negedge clk or negedge rst_n)
begin
   if(~rst_n)
      data_buf <= 8'd0;
   else if(start_bit_sig)
      data_buf <= din_byte;	 	           //din_byte;  // at just arriving the start_bit_sig , we load data into data_buffer 
   else if(data_bits_sig)
      data_buf <= {1'b1,data_buf[7:1]};
   else
      data_buf <= data_buf;
end
  
// Counter that count shift in Data Buffer Logic
always @(negedge clk or negedge rst_n)
begin
   if(~rst_n)
      shift_count <= 3'd0;
   else if(data_bits_sig)
      shift_count <= shift_count + 1; 
   else
      shift_count <= 3'd0;
end
// State machine for Tx
uat_sm uat_sm_inst(// Inputs
                   .clk              (clk),
                   .rst_n            (rst_n),
                   .din_rdy          (din_rdy_reg),      // 1-bit serial data from channel 
                   .shift_count      (shift_count),
                   // Outputs
                   .start_bit_sig    (start_bit_sig),    // Start bit insertion Control Signal generate from State Mechiene
                   .data_bits_sig    (data_bits_sig),    // Data bits insertion Control Signal generate from State Mechiene
                   .stop_bit_sig     (stop_bit_sig),     // Stop Bit insertion  Control Signal generate from State Mechiene
                   .uart_ready       (uart_ready) 
                  );
endmodule

